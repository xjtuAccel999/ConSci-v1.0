module LutZ
(
	input  logic [7:0]  index,
	output logic [24:0] lut_value
);

always_comb begin
    case (index)
		8'b00000000:	lut_value = 25'b0010110100010100001111110;
		8'b00000001:	lut_value = 25'b0010110011100111110001101;
		8'b00000010:	lut_value = 25'b0010110010111011110100001;
		8'b00000011:	lut_value = 25'b0010110010010000010110101;
		8'b00000100:	lut_value = 25'b0010110001100101011000100;
		8'b00000101:	lut_value = 25'b0010110000111010111001011;
		8'b00000110:	lut_value = 25'b0010110000010000111000100;
		8'b00000111:	lut_value = 25'b0010101111100111010101010;
		8'b00001000:	lut_value = 25'b0010101110111110001111001;
		8'b00001001:	lut_value = 25'b0010101110010101100101110;
		8'b00001010:	lut_value = 25'b0010101101101101011000100;
		8'b00001011:	lut_value = 25'b0010101101000101100110110;
		8'b00001100:	lut_value = 25'b0010101100011110010000010;
		8'b00001101:	lut_value = 25'b0010101011110111010100011;
		8'b00001110:	lut_value = 25'b0010101011010000110010101;
		8'b00001111:	lut_value = 25'b0010101010101010101010110;
		8'b00010000:	lut_value = 25'b0010101010000100111100000;
		8'b00010001:	lut_value = 25'b0010101001011111100110001;
		8'b00010010:	lut_value = 25'b0010101000111010101000110;
		8'b00010011:	lut_value = 25'b0010101000010110000011011;
		8'b00010100:	lut_value = 25'b0010100111110001110101100;
		8'b00010101:	lut_value = 25'b0010100111001101111111000;
		8'b00010110:	lut_value = 25'b0010100110101010011111010;
		8'b00010111:	lut_value = 25'b0010100110000111010101111;
		8'b00011000:	lut_value = 25'b0010100101100100100010110;
		8'b00011001:	lut_value = 25'b0010100101000010000101011;
		8'b00011010:	lut_value = 25'b0010100100011111111101010;
		8'b00011011:	lut_value = 25'b0010100011111110001010001;
		8'b00011100:	lut_value = 25'b0010100011011100101011110;
		8'b00011101:	lut_value = 25'b0010100010111011100001111;
		8'b00011110:	lut_value = 25'b0010100010011010101011111;
		8'b00011111:	lut_value = 25'b0010100001111010001001110;
		8'b00100000:	lut_value = 25'b0010100001011001111011000;
		8'b00100001:	lut_value = 25'b0010100000111001111111010;
		8'b00100010:	lut_value = 25'b0010100000011010010110100;
		8'b00100011:	lut_value = 25'b0010011111111011000000010;
		8'b00100100:	lut_value = 25'b0010011111011011111100010;
		8'b00100101:	lut_value = 25'b0010011110111101001010010;
		8'b00100110:	lut_value = 25'b0010011110011110101010000;
		8'b00100111:	lut_value = 25'b0010011110000000011011001;
		8'b00101000:	lut_value = 25'b0010011101100010011101100;
		8'b00101001:	lut_value = 25'b0010011101000100110000111;
		8'b00101010:	lut_value = 25'b0010011100100111010100111;
		8'b00101011:	lut_value = 25'b0010011100001010001001011;
		8'b00101100:	lut_value = 25'b0010011011101101001110001;
		8'b00101101:	lut_value = 25'b0010011011010000100010110;
		8'b00101110:	lut_value = 25'b0010011010110100000111001;
		8'b00101111:	lut_value = 25'b0010011010010111111011001;
		8'b00110000:	lut_value = 25'b0010011001111011111110011;
		8'b00110001:	lut_value = 25'b0010011001100000010000110;
		8'b00110010:	lut_value = 25'b0010011001000100110010000;
		8'b00110011:	lut_value = 25'b0010011000101001100001111;
		8'b00110100:	lut_value = 25'b0010011000001110100000010;
		8'b00110101:	lut_value = 25'b0010010111110011101101000;
		8'b00110110:	lut_value = 25'b0010010111011001000111110;
		8'b00110111:	lut_value = 25'b0010010110111110110000011;
		8'b00111000:	lut_value = 25'b0010010110100100100110110;
		8'b00111001:	lut_value = 25'b0010010110001010101010101;
		8'b00111010:	lut_value = 25'b0010010101110000111011110;
		8'b00111011:	lut_value = 25'b0010010101010111011010001;
		8'b00111100:	lut_value = 25'b0010010100111110000101100;
		8'b00111101:	lut_value = 25'b0010010100100100111101101;
		8'b00111110:	lut_value = 25'b0010010100001100000010011;
		8'b00111111:	lut_value = 25'b0010010011110011010011101;
		8'b01000000:	lut_value = 25'b0010010011011010110001010;
		8'b01000001:	lut_value = 25'b0010010011000010011011000;
		8'b01000010:	lut_value = 25'b0010010010101010010000110;
		8'b01000011:	lut_value = 25'b0010010010010010010010010;
		8'b01000100:	lut_value = 25'b0010010001111010011111100;
		8'b01000101:	lut_value = 25'b0010010001100010111000011;
		8'b01000110:	lut_value = 25'b0010010001001011011100101;
		8'b01000111:	lut_value = 25'b0010010000110100001100001;
		8'b01001000:	lut_value = 25'b0010010000011101000110110;
		8'b01001001:	lut_value = 25'b0010010000000110001100011;
		8'b01001010:	lut_value = 25'b0010001111101111011100111;
		8'b01001011:	lut_value = 25'b0010001111011000111000000;
		8'b01001100:	lut_value = 25'b0010001111000010011101110;
		8'b01001101:	lut_value = 25'b0010001110101100001110000;
		8'b01001110:	lut_value = 25'b0010001110010110001000100;
		8'b01001111:	lut_value = 25'b0010001110000000001101010;
		8'b01010000:	lut_value = 25'b0010001101101010011100001;
		8'b01010001:	lut_value = 25'b0010001101010100110101000;
		8'b01010010:	lut_value = 25'b0010001100111111010111101;
		8'b01010011:	lut_value = 25'b0010001100101010000100000;
		8'b01010100:	lut_value = 25'b0010001100010100111010000;
		8'b01010101:	lut_value = 25'b0010001011111111111001011;
		8'b01010110:	lut_value = 25'b0010001011101011000010010;
		8'b01010111:	lut_value = 25'b0010001011010110010100100;
		8'b01011000:	lut_value = 25'b0010001011000001101111111;
		8'b01011001:	lut_value = 25'b0010001010101101010100010;
		8'b01011010:	lut_value = 25'b0010001010011001000001101;
		8'b01011011:	lut_value = 25'b0010001010000100110111111;
		8'b01011100:	lut_value = 25'b0010001001110000110110111;
		8'b01011101:	lut_value = 25'b0010001001011100111110100;
		8'b01011110:	lut_value = 25'b0010001001001001001110110;
		8'b01011111:	lut_value = 25'b0010001000110101100111011;
		8'b01100000:	lut_value = 25'b0010001000100010001000100;
		8'b01100001:	lut_value = 25'b0010001000001110110001111;
		8'b01100010:	lut_value = 25'b0010000111111011100011100;
		8'b01100011:	lut_value = 25'b0010000111101000011101001;
		8'b01100100:	lut_value = 25'b0010000111010101011110110;
		8'b01100101:	lut_value = 25'b0010000111000010101000011;
		8'b01100110:	lut_value = 25'b0010000110101111111001111;
		8'b01100111:	lut_value = 25'b0010000110011101010011001;
		8'b01101000:	lut_value = 25'b0010000110001010110100000;
		8'b01101001:	lut_value = 25'b0010000101111000011100100;
		8'b01101010:	lut_value = 25'b0010000101100110001100100;
		8'b01101011:	lut_value = 25'b0010000101010100000011111;
		8'b01101100:	lut_value = 25'b0010000101000010000010101;
		8'b01101101:	lut_value = 25'b0010000100110000001000101;
		8'b01101110:	lut_value = 25'b0010000100011110010101111;
		8'b01101111:	lut_value = 25'b0010000100001100101010010;
		8'b01110000:	lut_value = 25'b0010000011111011000101110;
		8'b01110001:	lut_value = 25'b0010000011101001101000001;
		8'b01110010:	lut_value = 25'b0010000011011000010001011;
		8'b01110011:	lut_value = 25'b0010000011000111000001101;
		8'b01110100:	lut_value = 25'b0010000010110101111000100;
		8'b01110101:	lut_value = 25'b0010000010100100110110001;
		8'b01110110:	lut_value = 25'b0010000010010011111010011;
		8'b01110111:	lut_value = 25'b0010000010000011000101001;
		8'b01111000:	lut_value = 25'b0010000001110010010110011;
		8'b01111001:	lut_value = 25'b0010000001100001101110001;
		8'b01111010:	lut_value = 25'b0010000001010001001100010;
		8'b01111011:	lut_value = 25'b0010000001000000110000101;
		8'b01111100:	lut_value = 25'b0010000000110000011011010;
		8'b01111101:	lut_value = 25'b0010000000100000001100001;
		8'b01111110:	lut_value = 25'b0010000000010000000011000;
		8'b01111111:	lut_value = 25'b0010000000000000000000000;
		8'b10000000:	lut_value = 25'b0011111110000001011110111;
		8'b10000001:	lut_value = 25'b0011111110000001011110111;
		8'b10000010:	lut_value = 25'b0011111100000101110110011;
		8'b10000011:	lut_value = 25'b0011111100000101110110011;
		8'b10000100:	lut_value = 25'b0011111010001100111111101;
		8'b10000101:	lut_value = 25'b0011111010001100111111101;
		8'b10000110:	lut_value = 25'b0011111000010110110100001;
		8'b10000111:	lut_value = 25'b0011111000010110110100001;
		8'b10001000:	lut_value = 25'b0011110110100011001101110;
		8'b10001001:	lut_value = 25'b0011110110100011001101110;
		8'b10001010:	lut_value = 25'b0011110100110010000110011;
		8'b10001011:	lut_value = 25'b0011110100110010000110011;
		8'b10001100:	lut_value = 25'b0011110011000011011000101;
		8'b10001101:	lut_value = 25'b0011110011000011011000101;
		8'b10001110:	lut_value = 25'b0011110001010110111111000;
		8'b10001111:	lut_value = 25'b0011110001010110111111000;
		8'b10010000:	lut_value = 25'b0011101111101100110100010;
		8'b10010001:	lut_value = 25'b0011101111101100110100010;
		8'b10010010:	lut_value = 25'b0011101110000100110011111;
		8'b10010011:	lut_value = 25'b0011101110000100110011111;
		8'b10010100:	lut_value = 25'b0011101100011110111001000;
		8'b10010101:	lut_value = 25'b0011101100011110111001000;
		8'b10010110:	lut_value = 25'b0011101010111010111111011;
		8'b10010111:	lut_value = 25'b0011101010111010111111011;
		8'b10011000:	lut_value = 25'b0011101001011001000010101;
		8'b10011001:	lut_value = 25'b0011101001011001000010101;
		8'b10011010:	lut_value = 25'b0011100111111000111110111;
		8'b10011011:	lut_value = 25'b0011100111111000111110111;
		8'b10011100:	lut_value = 25'b0011100110011010110000001;
		8'b10011101:	lut_value = 25'b0011100110011010110000001;
		8'b10011110:	lut_value = 25'b0011100100111110010011000;
		8'b10011111:	lut_value = 25'b0011100100111110010011000;
		8'b10100000:	lut_value = 25'b0011100011100011100011100;
		8'b10100001:	lut_value = 25'b0011100011100011100011100;
		8'b10100010:	lut_value = 25'b0011100010001010011110110;
		8'b10100011:	lut_value = 25'b0011100010001010011110110;
		8'b10100100:	lut_value = 25'b0011100000110011000001011;
		8'b10100101:	lut_value = 25'b0011100000110011000001011;
		8'b10100110:	lut_value = 25'b0011011111011101001000010;
		8'b10100111:	lut_value = 25'b0011011111011101001000010;
		8'b10101000:	lut_value = 25'b0011011110001000110000010;
		8'b10101001:	lut_value = 25'b0011011110001000110000010;
		8'b10101010:	lut_value = 25'b0011011100110101110110111;
		8'b10101011:	lut_value = 25'b0011011100110101110110111;
		8'b10101100:	lut_value = 25'b0011011011100100011001010;
		8'b10101101:	lut_value = 25'b0011011011100100011001010;
		8'b10101110:	lut_value = 25'b0011011010010100010100101;
		8'b10101111:	lut_value = 25'b0011011010010100010100101;
		8'b10110000:	lut_value = 25'b0011011001000101100110101;
		8'b10110001:	lut_value = 25'b0011011001000101100110101;
		8'b10110010:	lut_value = 25'b0011010111111000001100111;
		8'b10110011:	lut_value = 25'b0011010111111000001100111;
		8'b10110100:	lut_value = 25'b0011010110101100000101001;
		8'b10110101:	lut_value = 25'b0011010110101100000101001;
		8'b10110110:	lut_value = 25'b0011010101100001001100111;
		8'b10110111:	lut_value = 25'b0011010101100001001100111;
		8'b10111000:	lut_value = 25'b0011010100010111100010001;
		8'b10111001:	lut_value = 25'b0011010100010111100010001;
		8'b10111010:	lut_value = 25'b0011010011001111000010111;
		8'b10111011:	lut_value = 25'b0011010011001111000010111;
		8'b10111100:	lut_value = 25'b0011010010000111101101000;
		8'b10111101:	lut_value = 25'b0011010010000111101101000;
		8'b10111110:	lut_value = 25'b0011010001000001011110110;
		8'b10111111:	lut_value = 25'b0011010001000001011110110;
		8'b11000000:	lut_value = 25'b0011001111111100010110000;
		8'b11000001:	lut_value = 25'b0011001111111100010110000;
		8'b11000010:	lut_value = 25'b0011001110111000010001011;
		8'b11000011:	lut_value = 25'b0011001110111000010001011;
		8'b11000100:	lut_value = 25'b0011001101110101001110111;
		8'b11000101:	lut_value = 25'b0011001101110101001110111;
		8'b11000110:	lut_value = 25'b0011001100110011001100110;
		8'b11000111:	lut_value = 25'b0011001100110011001100110;
		8'b11001000:	lut_value = 25'b0011001011110010001001110;
		8'b11001001:	lut_value = 25'b0011001011110010001001110;
		8'b11001010:	lut_value = 25'b0011001010110010000100000;
		8'b11001011:	lut_value = 25'b0011001010110010000100000;
		8'b11001100:	lut_value = 25'b0011001001110010111010001;
		8'b11001101:	lut_value = 25'b0011001001110010111010001;
		8'b11001110:	lut_value = 25'b0011001000110100101010101;
		8'b11001111:	lut_value = 25'b0011001000110100101010101;
		8'b11010000:	lut_value = 25'b0011000111110111010100011;
		8'b11010001:	lut_value = 25'b0011000111110111010100011;
		8'b11010010:	lut_value = 25'b0011000110111010110101101;
		8'b11010011:	lut_value = 25'b0011000110111010110101101;
		8'b11010100:	lut_value = 25'b0011000101111111001101011;
		8'b11010101:	lut_value = 25'b0011000101111111001101011;
		8'b11010110:	lut_value = 25'b0011000101000100011010001;
		8'b11010111:	lut_value = 25'b0011000101000100011010001;
		8'b11011000:	lut_value = 25'b0011000100001010011011000;
		8'b11011001:	lut_value = 25'b0011000100001010011011000;
		8'b11011010:	lut_value = 25'b0011000011010001001110011;
		8'b11011011:	lut_value = 25'b0011000011010001001110011;
		8'b11011100:	lut_value = 25'b0011000010011000110011100;
		8'b11011101:	lut_value = 25'b0011000010011000110011100;
		8'b11011110:	lut_value = 25'b0011000001100001001001000;
		8'b11011111:	lut_value = 25'b0011000001100001001001000;
		8'b11100000:	lut_value = 25'b0011000000101010001101111;
		8'b11100001:	lut_value = 25'b0011000000101010001101111;
		8'b11100010:	lut_value = 25'b0010111111110100000001001;
		8'b11100011:	lut_value = 25'b0010111111110100000001001;
		8'b11100100:	lut_value = 25'b0010111110111110100001110;
		8'b11100101:	lut_value = 25'b0010111110111110100001110;
		8'b11100110:	lut_value = 25'b0010111110001001101110101;
		8'b11100111:	lut_value = 25'b0010111110001001101110101;
		8'b11101000:	lut_value = 25'b0010111101010101100111001;
		8'b11101001:	lut_value = 25'b0010111101010101100111001;
		8'b11101010:	lut_value = 25'b0010111100100010001001111;
		8'b11101011:	lut_value = 25'b0010111100100010001001111;
		8'b11101100:	lut_value = 25'b0010111011101111010110100;
		8'b11101101:	lut_value = 25'b0010111011101111010110100;
		8'b11101110:	lut_value = 25'b0010111010111101001011101;
		8'b11101111:	lut_value = 25'b0010111010111101001011101;
		8'b11110000:	lut_value = 25'b0010111010001011101000110;
		8'b11110001:	lut_value = 25'b0010111010001011101000110;
		8'b11110010:	lut_value = 25'b0010111001011010101100111;
		8'b11110011:	lut_value = 25'b0010111001011010101100111;
		8'b11110100:	lut_value = 25'b0010111000101010010111010;
		8'b11110101:	lut_value = 25'b0010111000101010010111010;
		8'b11110110:	lut_value = 25'b0010110111111010100111010;
		8'b11110111:	lut_value = 25'b0010110111111010100111010;
		8'b11111000:	lut_value = 25'b0010110111001011011011111;
		8'b11111001:	lut_value = 25'b0010110111001011011011111;
		8'b11111010:	lut_value = 25'b0010110110011100110100101;
		8'b11111011:	lut_value = 25'b0010110110011100110100101;
		8'b11111100:	lut_value = 25'b0010110101101110110000101;
		8'b11111101:	lut_value = 25'b0010110101101110110000101;
		8'b11111110:	lut_value = 25'b0010110101000001001111001;
		8'b11111111:	lut_value = 25'b0010110101000001001111001;
	endcase
end
endmodule

module LutZ3
(
	input  logic [7:0]  index,
	output logic [24:0] lut_value
);

always_comb begin
    case (index)
		8'b00000000:	lut_value = 25'b0001011001011101011001000;
		8'b00000001:	lut_value = 25'b0001011000011011011101010;
		8'b00000010:	lut_value = 25'b0001010111011010110001110;
		8'b00000011:	lut_value = 25'b0001010110011011010100101;
		8'b00000100:	lut_value = 25'b0001010101011101000011011;
		8'b00000101:	lut_value = 25'b0001010100011111111100110;
		8'b00000110:	lut_value = 25'b0001010011100011111110011;
		8'b00000111:	lut_value = 25'b0001010010101001000110001;
		8'b00001000:	lut_value = 25'b0001010001101111010010101;
		8'b00001001:	lut_value = 25'b0001010000110110100010001;
		8'b00001010:	lut_value = 25'b0001001111111110110010111;
		8'b00001011:	lut_value = 25'b0001001111001000000010111;
		8'b00001100:	lut_value = 25'b0001001110010010010001010;
		8'b00001101:	lut_value = 25'b0001001101011101011100000;
		8'b00001110:	lut_value = 25'b0001001100101001100001110;
		8'b00001111:	lut_value = 25'b0001001011110110100001010;
		8'b00010000:	lut_value = 25'b0001001011000100011000101;
		8'b00010001:	lut_value = 25'b0001001010010011000110111;
		8'b00010010:	lut_value = 25'b0001001001100010101010111;
		8'b00010011:	lut_value = 25'b0001001000110011000011001;
		8'b00010100:	lut_value = 25'b0001001000000100001110010;
		8'b00010101:	lut_value = 25'b0001000111010110001011011;
		8'b00010110:	lut_value = 25'b0001000110101000111001010;
		8'b00010111:	lut_value = 25'b0001000101111100010110100;
		8'b00011000:	lut_value = 25'b0001000101010000100010100;
		8'b00011001:	lut_value = 25'b0001000100100101011100000;
		8'b00011010:	lut_value = 25'b0001000011111011000001101;
		8'b00011011:	lut_value = 25'b0001000011010001010010110;
		8'b00011100:	lut_value = 25'b0001000010101000001110011;
		8'b00011101:	lut_value = 25'b0001000001111111110011110;
		8'b00011110:	lut_value = 25'b0001000001011000000001100;
		8'b00011111:	lut_value = 25'b0001000000110000110111000;
		8'b00100000:	lut_value = 25'b0001000000001010010011011;
		8'b00100001:	lut_value = 25'b0000111111100100010101110;
		8'b00100010:	lut_value = 25'b0000111110111110111101011;
		8'b00100011:	lut_value = 25'b0000111110011010001001011;
		8'b00100100:	lut_value = 25'b0000111101110101111001000;
		8'b00100101:	lut_value = 25'b0000111101010010001011101;
		8'b00100110:	lut_value = 25'b0000111100101111000000011;
		8'b00100111:	lut_value = 25'b0000111100001100010110011;
		8'b00101000:	lut_value = 25'b0000111011101010001101010;
		8'b00101001:	lut_value = 25'b0000111011001000100100011;
		8'b00101010:	lut_value = 25'b0000111010100111011010110;
		8'b00101011:	lut_value = 25'b0000111010000110110000000;
		8'b00101100:	lut_value = 25'b0000111001100110100011100;
		8'b00101101:	lut_value = 25'b0000111001000110110100100;
		8'b00101110:	lut_value = 25'b0000111000100111100010010;
		8'b00101111:	lut_value = 25'b0000111000001000101100101;
		8'b00110000:	lut_value = 25'b0000110111101010010010110;
		8'b00110001:	lut_value = 25'b0000110111001100010100010;
		8'b00110010:	lut_value = 25'b0000110110101110110000100;
		8'b00110011:	lut_value = 25'b0000110110010001100110111;
		8'b00110100:	lut_value = 25'b0000110101110100110111001;
		8'b00110101:	lut_value = 25'b0000110101011000100000101;
		8'b00110110:	lut_value = 25'b0000110100111100100010110;
		8'b00110111:	lut_value = 25'b0000110100100000111101010;
		8'b00111000:	lut_value = 25'b0000110100000101101111101;
		8'b00111001:	lut_value = 25'b0000110011101010111001010;
		8'b00111010:	lut_value = 25'b0000110011010000011001111;
		8'b00111011:	lut_value = 25'b0000110010110110010001000;
		8'b00111100:	lut_value = 25'b0000110010011100011110010;
		8'b00111101:	lut_value = 25'b0000110010000011000001001;
		8'b00111110:	lut_value = 25'b0000110001101001111001011;
		8'b00111111:	lut_value = 25'b0000110001010001000110011;
		8'b01000000:	lut_value = 25'b0000110000111000101000001;
		8'b01000001:	lut_value = 25'b0000110000100000011110000;
		8'b01000010:	lut_value = 25'b0000110000001000100111100;
		8'b01000011:	lut_value = 25'b0000101111110001000100100;
		8'b01000100:	lut_value = 25'b0000101111011001110100101;
		8'b01000101:	lut_value = 25'b0000101111000010110111101;
		8'b01000110:	lut_value = 25'b0000101110101100001101000;
		8'b01000111:	lut_value = 25'b0000101110010101110100011;
		8'b01001000:	lut_value = 25'b0000101101111111101101101;
		8'b01001001:	lut_value = 25'b0000101101101001111000011;
		8'b01001010:	lut_value = 25'b0000101101010100010100011;
		8'b01001011:	lut_value = 25'b0000101100111111000001001;
		8'b01001100:	lut_value = 25'b0000101100101001111110101;
		8'b01001101:	lut_value = 25'b0000101100010101001100011;
		8'b01001110:	lut_value = 25'b0000101100000000101010000;
		8'b01001111:	lut_value = 25'b0000101011101100010111101;
		8'b01010000:	lut_value = 25'b0000101011011000010100110;
		8'b01010001:	lut_value = 25'b0000101011000100100001001;
		8'b01010010:	lut_value = 25'b0000101010110000111100100;
		8'b01010011:	lut_value = 25'b0000101010011101100110101;
		8'b01010100:	lut_value = 25'b0000101010001010011111010;
		8'b01010101:	lut_value = 25'b0000101001110111100110000;
		8'b01010110:	lut_value = 25'b0000101001100100111010111;
		8'b01010111:	lut_value = 25'b0000101001010010011101101;
		8'b01011000:	lut_value = 25'b0000101001000000001110001;
		8'b01011001:	lut_value = 25'b0000101000101110001011110;
		8'b01011010:	lut_value = 25'b0000101000011100010110101;
		8'b01011011:	lut_value = 25'b0000101000001010101110011;
		8'b01011100:	lut_value = 25'b0000100111111001010011000;
		8'b01011101:	lut_value = 25'b0000100111101000000100001;
		8'b01011110:	lut_value = 25'b0000100111010111000001100;
		8'b01011111:	lut_value = 25'b0000100111000110001011001;
		8'b01100000:	lut_value = 25'b0000100110110101100000110;
		8'b01100001:	lut_value = 25'b0000100110100101000010001;
		8'b01100010:	lut_value = 25'b0000100110010100101111001;
		8'b01100011:	lut_value = 25'b0000100110000100100111100;
		8'b01100100:	lut_value = 25'b0000100101110100101011001;
		8'b01100101:	lut_value = 25'b0000100101100100111001111;
		8'b01100110:	lut_value = 25'b0000100101010101010011100;
		8'b01100111:	lut_value = 25'b0000100101000101110111111;
		8'b01101000:	lut_value = 25'b0000100100110110100111000;
		8'b01101001:	lut_value = 25'b0000100100100111100000011;
		8'b01101010:	lut_value = 25'b0000100100011000100100000;
		8'b01101011:	lut_value = 25'b0000100100001001110001110;
		8'b01101100:	lut_value = 25'b0000100011111011001001100;
		8'b01101101:	lut_value = 25'b0000100011101100101011000;
		8'b01101110:	lut_value = 25'b0000100011011110010110011;
		8'b01101111:	lut_value = 25'b0000100011010000001011001;
		8'b01110000:	lut_value = 25'b0000100011000010001001011;
		8'b01110001:	lut_value = 25'b0000100010110100010000111;
		8'b01110010:	lut_value = 25'b0000100010100110100001011;
		8'b01110011:	lut_value = 25'b0000100010011000111011001;
		8'b01110100:	lut_value = 25'b0000100010001011011101100;
		8'b01110101:	lut_value = 25'b0000100001111110001000110;
		8'b01110110:	lut_value = 25'b0000100001110000111100101;
		8'b01110111:	lut_value = 25'b0000100001100011111000111;
		8'b01111000:	lut_value = 25'b0000100001010110111101101;
		8'b01111001:	lut_value = 25'b0000100001001010001010101;
		8'b01111010:	lut_value = 25'b0000100000111101011111111;
		8'b01111011:	lut_value = 25'b0000100000110000111101000;
		8'b01111100:	lut_value = 25'b0000100000100100100010001;
		8'b01111101:	lut_value = 25'b0000100000011000001111001;
		8'b01111110:	lut_value = 25'b0000100000001100000011110;
		8'b01111111:	lut_value = 25'b0000100000000000000000000;
		8'b10000000:	lut_value = 25'b0011111010000111010111101;
		8'b10000001:	lut_value = 25'b0011111010000111010111101;
		8'b10000010:	lut_value = 25'b0011110100011100111100101;
		8'b10000011:	lut_value = 25'b0011110100011100111100101;
		8'b10000100:	lut_value = 25'b0011101110111111111111101;
		8'b10000101:	lut_value = 25'b0011101110111111111111101;
		8'b10000110:	lut_value = 25'b0011101001101111110100110;
		8'b10000111:	lut_value = 25'b0011101001101111110100110;
		8'b10001000:	lut_value = 25'b0011100100101011110010110;
		8'b10001001:	lut_value = 25'b0011100100101011110010110;
		8'b10001010:	lut_value = 25'b0011011111110011010010011;
		8'b10001011:	lut_value = 25'b0011011111110011010010011;
		8'b10001100:	lut_value = 25'b0011011011000101110000010;
		8'b10001101:	lut_value = 25'b0011011011000101110000010;
		8'b10001110:	lut_value = 25'b0011010110100010101001110;
		8'b10001111:	lut_value = 25'b0011010110100010101001110;
		8'b10010000:	lut_value = 25'b0011010010001001011110110;
		8'b10010001:	lut_value = 25'b0011010010001001011110110;
		8'b10010010:	lut_value = 25'b0011001101111001110010000;
		8'b10010011:	lut_value = 25'b0011001101111001110010000;
		8'b10010100:	lut_value = 25'b0011001001110011000110101;
		8'b10010101:	lut_value = 25'b0011001001110011000110101;
		8'b10010110:	lut_value = 25'b0011000101110101000010110;
		8'b10010111:	lut_value = 25'b0011000101110101000010110;
		8'b10011000:	lut_value = 25'b0011000001111111001100111;
		8'b10011001:	lut_value = 25'b0011000001111111001100111;
		8'b10011010:	lut_value = 25'b0010111110010001001101111;
		8'b10011011:	lut_value = 25'b0010111110010001001101111;
		8'b10011100:	lut_value = 25'b0010111010101010101111000;
		8'b10011101:	lut_value = 25'b0010111010101010101111000;
		8'b10011110:	lut_value = 25'b0010110111001011011100001;
		8'b10011111:	lut_value = 25'b0010110111001011011100001;
		8'b10100000:	lut_value = 25'b0010110011110011000000010;
		8'b10100001:	lut_value = 25'b0010110011110011000000010;
		8'b10100010:	lut_value = 25'b0010110000100001001001110;
		8'b10100011:	lut_value = 25'b0010110000100001001001110;
		8'b10100100:	lut_value = 25'b0010101101010101100110110;
		8'b10100101:	lut_value = 25'b0010101101010101100110110;
		8'b10100110:	lut_value = 25'b0010101010010000000110010;
		8'b10100111:	lut_value = 25'b0010101010010000000110010;
		8'b10101000:	lut_value = 25'b0010100111010000011000001;
		8'b10101001:	lut_value = 25'b0010100111010000011000001;
		8'b10101010:	lut_value = 25'b0010100100010110001110000;
		8'b10101011:	lut_value = 25'b0010100100010110001110000;
		8'b10101100:	lut_value = 25'b0010100001100001011001010;
		8'b10101101:	lut_value = 25'b0010100001100001011001010;
		8'b10101110:	lut_value = 25'b0010011110110001101100000;
		8'b10101111:	lut_value = 25'b0010011110110001101100000;
		8'b10110000:	lut_value = 25'b0010011100000110111001110;
		8'b10110001:	lut_value = 25'b0010011100000110111001110;
		8'b10110010:	lut_value = 25'b0010011001100000110110100;
		8'b10110011:	lut_value = 25'b0010011001100000110110100;
		8'b10110100:	lut_value = 25'b0010010110111111010110101;
		8'b10110101:	lut_value = 25'b0010010110111111010110101;
		8'b10110110:	lut_value = 25'b0010010100100010001110011;
		8'b10110111:	lut_value = 25'b0010010100100010001110011;
		8'b10111000:	lut_value = 25'b0010010010001001010011111;
		8'b10111001:	lut_value = 25'b0010010010001001010011111;
		8'b10111010:	lut_value = 25'b0010001111110100011101000;
		8'b10111011:	lut_value = 25'b0010001111110100011101000;
		8'b10111100:	lut_value = 25'b0010001101100011100000010;
		8'b10111101:	lut_value = 25'b0010001101100011100000010;
		8'b10111110:	lut_value = 25'b0010001011010110010100011;
		8'b10111111:	lut_value = 25'b0010001011010110010100011;
		8'b11000000:	lut_value = 25'b0010001001001100110000101;
		8'b11000001:	lut_value = 25'b0010001001001100110000101;
		8'b11000010:	lut_value = 25'b0010000111000110101101001;
		8'b11000011:	lut_value = 25'b0010000111000110101101001;
		8'b11000100:	lut_value = 25'b0010000101000100000001111;
		8'b11000101:	lut_value = 25'b0010000101000100000001111;
		8'b11000110:	lut_value = 25'b0010000011000100100110110;
		8'b11000111:	lut_value = 25'b0010000011000100100110110;
		8'b11001000:	lut_value = 25'b0010000001001000010101011;
		8'b11001001:	lut_value = 25'b0010000001001000010101011;
		8'b11001010:	lut_value = 25'b0001111111001111000110001;
		8'b11001011:	lut_value = 25'b0001111111001111000110001;
		8'b11001100:	lut_value = 25'b0001111101011000110011000;
		8'b11001101:	lut_value = 25'b0001111101011000110011000;
		8'b11001110:	lut_value = 25'b0001111011100101010101001;
		8'b11001111:	lut_value = 25'b0001111011100101010101001;
		8'b11010000:	lut_value = 25'b0001111001110100100111010;
		8'b11010001:	lut_value = 25'b0001111001110100100111010;
		8'b11010010:	lut_value = 25'b0001111000000110100010101;
		8'b11010011:	lut_value = 25'b0001111000000110100010101;
		8'b11010100:	lut_value = 25'b0001110110011011000010100;
		8'b11010101:	lut_value = 25'b0001110110011011000010100;
		8'b11010110:	lut_value = 25'b0001110100110010000001001;
		8'b11010111:	lut_value = 25'b0001110100110010000001001;
		8'b11011000:	lut_value = 25'b0001110011001011011001111;
		8'b11011001:	lut_value = 25'b0001110011001011011001111;
		8'b11011010:	lut_value = 25'b0001110001100111000111001;
		8'b11011011:	lut_value = 25'b0001110001100111000111001;
		8'b11011100:	lut_value = 25'b0001110000000101000100111;
		8'b11011101:	lut_value = 25'b0001110000000101000100111;
		8'b11011110:	lut_value = 25'b0001101110100101001110010;
		8'b11011111:	lut_value = 25'b0001101110100101001110010;
		8'b11100000:	lut_value = 25'b0001101101000111011111000;
		8'b11100001:	lut_value = 25'b0001101101000111011111000;
		8'b11100010:	lut_value = 25'b0001101011101011110011000;
		8'b11100011:	lut_value = 25'b0001101011101011110011000;
		8'b11100100:	lut_value = 25'b0001101010010010000110011;
		8'b11100101:	lut_value = 25'b0001101010010010000110011;
		8'b11100110:	lut_value = 25'b0001101000111010010101001;
		8'b11100111:	lut_value = 25'b0001101000111010010101001;
		8'b11101000:	lut_value = 25'b0001100111100100011011111;
		8'b11101001:	lut_value = 25'b0001100111100100011011111;
		8'b11101010:	lut_value = 25'b0001100110010000010110100;
		8'b11101011:	lut_value = 25'b0001100110010000010110100;
		8'b11101100:	lut_value = 25'b0001100100111110000010011;
		8'b11101101:	lut_value = 25'b0001100100111110000010011;
		8'b11101110:	lut_value = 25'b0001100011101101011011100;
		8'b11101111:	lut_value = 25'b0001100011101101011011100;
		8'b11110000:	lut_value = 25'b0001100010011110011111000;
		8'b11110001:	lut_value = 25'b0001100010011110011111000;
		8'b11110010:	lut_value = 25'b0001100001010001001001111;
		8'b11110011:	lut_value = 25'b0001100001010001001001111;
		8'b11110100:	lut_value = 25'b0001100000000101011001000;
		8'b11110101:	lut_value = 25'b0001100000000101011001000;
		8'b11110110:	lut_value = 25'b0001011110111011001001111;
		8'b11110111:	lut_value = 25'b0001011110111011001001111;
		8'b11111000:	lut_value = 25'b0001011101110010011001011;
		8'b11111001:	lut_value = 25'b0001011101110010011001011;
		8'b11111010:	lut_value = 25'b0001011100101011000101010;
		8'b11111011:	lut_value = 25'b0001011100101011000101010;
		8'b11111100:	lut_value = 25'b0001011011100101001010111;
		8'b11111101:	lut_value = 25'b0001011011100101001010111;
		8'b11111110:	lut_value = 25'b0001011010100000100111011;
		8'b11111111:	lut_value = 25'b0001011010100000100111011;
	endcase
end
endmodule

module math_sqrtf32
(
	input logic 		clk,
	input logic 		rst_n,
	input logic 		sqrt_op_en,
	input logic [31:0] 	sqrt_rb,
	output logic 		sqrt_ra_en,
	output logic [31:0] sqrt_ra,
	output logic 		sqrt_lvf_flag
);

/* shift reg for pipeline */
logic [4:0] shift_reg_sqrt;

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n)
		shift_reg_sqrt <= 5'b0;
	else
		shift_reg_sqrt <= {shift_reg_sqrt[3:0], sqrt_op_en};
end

// Pipeline Level 1
/* Process Exponent */
logic [7:0] exp;
assign exp = sqrt_rb[23] ? sqrt_rb[30:24] + 8'd64 : sqrt_rb[30:24] + 8'd63;

/* Preprocess Tail */
logic [31:0] enabled_sqrt_rb;
logic [7:0] index;
logic [24:0] B;
logic [24:0] Z;
logic [24:0] Z3;
logic [55:0] BZ3;
logic [27:0] temp_x;
logic [27:0] temp_x1;

logic minus_flag;
logic inf_flag;
logic zero_flag;

assign enabled_sqrt_rb = sqrt_op_en ? sqrt_rb : 32'h00000000;
assign minus_flag 	= enabled_sqrt_rb[31];
assign inf_flag 	= (enabled_sqrt_rb[30:23] == 8'hff) ? 1'b1 : 1'b0;
assign zero_flag 	= (enabled_sqrt_rb[30:23] == 8'h00) ? 1'b1 : 1'b0;

assign index = enabled_sqrt_rb[23:16];
assign B = enabled_sqrt_rb[23] ? {2'b01, enabled_sqrt_rb[22:0]} : {1'b1, enabled_sqrt_rb[22:0], 1'b0};

LutZ u_LutZ
(
	.index		(	index		),
	.lut_value	(	Z			)
);

LutZ3 u_LutZ3
(
	.index		(	index		),
	.lut_value	(	Z3			)
);


assign BZ3 		= {B, 3'b0} * {Z3, 3'b0};
assign temp_x 	= {Z, 3'b0} + {Z[23:0], 4'b0} - BZ3[53:26];
assign temp_x1 	= {1'b0, temp_x[27:1]};

//Pipeline Register
logic [27:0] reg_X1_L1;
logic [24:0] reg_B_L1;
logic [7:0] reg_exp_L1;
logic reg_minus_flag_L1; 
logic reg_inf_flag_L1;
logic reg_zero_flag_L1;

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n) begin
		reg_X1_L1	<=	28'h0;
		reg_B_L1	<=	25'h0;	
		reg_exp_L1	<=	8'h0;
		reg_minus_flag_L1	<=	1'h0; 
		reg_inf_flag_L1		<=	1'h0;
		reg_zero_flag_L1	<=	1'h0;
	end
	else begin
		reg_X1_L1	<=	temp_x1;
		reg_B_L1	<=	B;
		reg_exp_L1	<=	exp;
		reg_minus_flag_L1	<=	minus_flag; 
		reg_inf_flag_L1		<=	inf_flag;
		reg_zero_flag_L1	<=	zero_flag;
	end
end	

// Pipeline Level 2
logic [55:0] temp_y1;

logic [27:0] reg_X1_L2;
logic [24:0] reg_B_L2;
logic [27:0] reg_Y1_L2;
logic [7:0] reg_exp_L2;
logic reg_minus_flag_L2; 
logic reg_inf_flag_L2;
logic reg_zero_flag_L2;

assign temp_y1 = reg_X1_L1 * {reg_B_L1, 3'b0};

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n) begin
		reg_X1_L2	<=	28'h0;
		reg_B_L2	<=	25'h0;
		reg_Y1_L2	<=	28'h0;
		reg_exp_L2	<=	8'h0;
		reg_minus_flag_L2	<= 1'h0; 
		reg_inf_flag_L2		<= 1'h0;
		reg_zero_flag_L2	<= 1'h0;
	end
	else begin
		reg_X1_L2	<=	reg_X1_L1;
		reg_B_L2	<=	reg_B_L1;
		reg_Y1_L2	<=	temp_y1[53:26];
		reg_exp_L2	<=	reg_exp_L1;
		reg_minus_flag_L2	<= reg_minus_flag_L1; 
		reg_inf_flag_L2		<= reg_inf_flag_L1;
		reg_zero_flag_L2	<= reg_zero_flag_L1;
	end
end	

// Pipeline Level 3
logic [55:0] temp_xy;
logic [27:0] temp_sub;

logic [27:0] reg_T0_L3;
logic [27:0] reg_Y1_L3;
logic [24:0] reg_B_L3;
logic [7:0]  reg_exp_L3;
logic reg_minus_flag_L3; 
logic reg_inf_flag_L3;
logic reg_zero_flag_L3;

parameter THREE = 28'b1100000000000000000000000000;

assign temp_xy = reg_X1_L2 * reg_Y1_L2;
assign temp_sub = THREE - temp_xy[53:26];

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n) begin
		reg_T0_L3	<= 28'h0;
		reg_Y1_L3	<= 28'h0;
		reg_B_L3	<= 25'h0;
		reg_exp_L3	<= 8'h0;
		reg_minus_flag_L3	<= 1'h0; 
		reg_inf_flag_L3		<= 1'h0;
		reg_zero_flag_L3	<= 1'h0;
	end 
	else begin 
		reg_T0_L3	<= temp_sub;
		reg_Y1_L3	<= reg_Y1_L2;
		reg_B_L3	<= reg_B_L2;
		reg_exp_L3	<= reg_exp_L2;	
		reg_minus_flag_L3	<= reg_minus_flag_L2; 
		reg_inf_flag_L3		<= reg_inf_flag_L2;
		reg_zero_flag_L3	<= reg_zero_flag_L2;
	end
end

// Pipeline Level 4
logic [55:0] temp_yt;
logic [27:0] temp_t;

logic [27:0] reg_T_L4;
logic [24:0] reg_B_L4;
logic [7:0]  reg_exp_L4;
logic reg_minus_flag_L4; 
logic reg_inf_flag_L4;
logic reg_zero_flag_L4;

logic temp_overflow_flag;
logic overflow_flag;

assign temp_yt = reg_T0_L3 * reg_Y1_L3;
assign temp_t = {1'b0, temp_yt[53:27]};

assign temp_overflow_flag = (reg_minus_flag_L3 | reg_inf_flag_L3) & ~reg_zero_flag_L3;

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n)
		overflow_flag <= 1'b0;
	else
		overflow_flag <= temp_overflow_flag;
end

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n) begin
		reg_T_L4	<= 28'h0;
		reg_B_L4	<= 25'h0;
		reg_exp_L4	<= 8'h0;
		reg_minus_flag_L4	<= 1'h0; 
		reg_inf_flag_L4		<= 1'h0;
		reg_zero_flag_L4	<= 1'h0;
	end 
	else begin 
		reg_T_L4	<= temp_t;
		reg_B_L4	<= reg_B_L3;
		reg_exp_L4	<= reg_exp_L3;	
		reg_minus_flag_L4	<= reg_minus_flag_L3; 
		reg_inf_flag_L4		<= reg_inf_flag_L3;
		reg_zero_flag_L4	<= reg_zero_flag_L3;
	end
end

// Pipeline Level 5
logic [24:0] R;
logic [49:0] R_square;
logic [50:0] D1, D2;
logic [24:0] R_plus_1;
logic [24:0] R_minus_1;
logic bor1, bor2;

logic [24:0] R_new;
logic [7:0] ra_exp;
logic [22:0] ra_tail;

logic [31:0] output_value;

assign R 		 = reg_T_L4[27:3];
assign R_square  = R * R;
assign R_plus_1  = R + 1'b1;
assign R_minus_1 = R - 1'b1;
assign D1		 = {reg_B_L4, 23'b0} + R - R_square;
assign D2		 = R_square + R - {reg_B_L4, 23'b0};
assign bor1		 = D1[50];
assign bor2		 = D2[50];

always_comb begin
	case({bor1, bor2})
		2'b00:		R_new = R;
		2'b01:		R_new = R_plus_1;
		2'b10:		R_new = R_minus_1;
		2'b11:		R_new = R;
		default:	R_new = R;
	endcase	
end

always_comb begin
	if (reg_zero_flag_L4)
		ra_exp = 8'h00;
	else if (reg_minus_flag_L4)
		ra_exp = 8'h00;
	else if (reg_inf_flag_L4)
		ra_exp = 8'hff;
	else
		ra_exp = reg_exp_L4;
end

always_comb begin
	if (reg_zero_flag_L4)
		ra_tail = 23'h0;
	else if (reg_minus_flag_L4)
		ra_tail = 23'h0;
	else if (reg_inf_flag_L4)
		ra_tail = 23'h0;
	else
		ra_tail = R_new;
end		

always_ff @(posedge clk or negedge rst_n)
begin
	if (~rst_n)
		output_value <= 32'h0;
	else if (shift_reg_sqrt[3])
		output_value <= {1'b0, ra_exp, ra_tail};
	else
		output_value <= output_value;
end

assign sqrt_ra 		 = 	output_value;
assign sqrt_ra_en	 =	shift_reg_sqrt[4];
assign sqrt_lvf_flag =	overflow_flag;
endmodule
