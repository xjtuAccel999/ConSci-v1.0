module mult_exp(
	input wire [31:0] mult_a,
	input wire [31:0] mult_b,
	output wire [31:0] mult_c
);

	wire [63:0] mult_temp;
	assign mult_temp = mult_a * mult_b;
	assign mult_c = mult_temp[63] ? mult_temp[63:32] : mult_temp[62:31];
endmodule  

module Lut1_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111101001111100000110000001100;
		6'b000010: lut_value = 32'b11111010100000111011001011011011;
		6'b000011: lut_value = 32'b11110111110100001101111101110011;
		6'b000100: lut_value = 32'b11110101001001010111110100010101;
		6'b000101: lut_value = 32'b11110010100000010111011100111100;
		6'b000110: lut_value = 32'b11101111111001001011100110011011;
		6'b000111: lut_value = 32'b11101101010011110011000000011110;
		6'b001000: lut_value = 32'b11101010110000001100011011100111;
		6'b001001: lut_value = 32'b11101000001110010110101001010000;
		6'b001010: lut_value = 32'b11100101101110010000011011100111;
		6'b001011: lut_value = 32'b11100011001111111000100101110010;
		6'b001100: lut_value = 32'b11100000110011001101111011101100;
		6'b001101: lut_value = 32'b11011110011000001111010010000010;
		6'b001110: lut_value = 32'b11011011111110111011011110010111;
		6'b001111: lut_value = 32'b11011001100111010001010111000010;
		6'b010000: lut_value = 32'b11010111010001001111110011001010;
		6'b010001: lut_value = 32'b11010100111100110101101010101011;
		6'b010010: lut_value = 32'b11010010101010000001110110010001;
		6'b010011: lut_value = 32'b11010000011000110011001111011010;
		6'b010100: lut_value = 32'b11001110001001001000110000010101;
		6'b010101: lut_value = 32'b11001011111011000001010011111110;
		6'b010110: lut_value = 32'b11001001101110011011110110000110;
		6'b010111: lut_value = 32'b11000111100011010111010011001000;
		6'b011000: lut_value = 32'b11000101011001110010101000010001;
		6'b011001: lut_value = 32'b11000011010001101100110011011010;
		6'b011010: lut_value = 32'b11000001001011000100110011001010;
		6'b011011: lut_value = 32'b10111111000101111001100110110110;
		6'b011100: lut_value = 32'b10111101000010001010001110011111;
		6'b011101: lut_value = 32'b10111010111111110101101010110010;
		6'b011110: lut_value = 32'b10111000111110111010111101000111;
		6'b011111: lut_value = 32'b10110110111111011001000111100011;
		6'b100000: lut_value = 32'b10110101000001001111001100110011;
		6'b100001: lut_value = 32'b10110011000100011100010000010010;
		6'b100010: lut_value = 32'b10110001001000111111010110000001;
		6'b100011: lut_value = 32'b10101111001110110111100010101101;
		6'b100100: lut_value = 32'b10101101010110000011111011101010;
		6'b100101: lut_value = 32'b10101011011110100011100110110101;
		6'b100110: lut_value = 32'b10101001101000010101101010110100;
		6'b100111: lut_value = 32'b10100111110011011001001110110100;
		6'b101000: lut_value = 32'b10100101111111101101011010101001;
		6'b101001: lut_value = 32'b10100100001101010001010110101110;
		6'b101010: lut_value = 32'b10100010011100000100001100000011;
		6'b101011: lut_value = 32'b10100000101100000101000100001111;
		6'b101100: lut_value = 32'b10011110111101010011001001100000;
		6'b101101: lut_value = 32'b10011101001111101101100110100111;
		6'b101110: lut_value = 32'b10011011100011010011100110111001;
		6'b101111: lut_value = 32'b10011001111000000100010110010011;
		6'b110000: lut_value = 32'b10011000001101111111000001010001;
		6'b110001: lut_value = 32'b10010110100101000010110100110111;
		6'b110010: lut_value = 32'b10010100111101001110111110101000;
		6'b110011: lut_value = 32'b10010011010110100010101100101111;
		6'b110100: lut_value = 32'b10010001110000111101001101110011;
		6'b110101: lut_value = 32'b10010000001100011101110001000011;
		6'b110110: lut_value = 32'b10001110101001000011100110001011;
		6'b110111: lut_value = 32'b10001101000110101101111101011011;
		6'b111000: lut_value = 32'b10001011100101011100000111100011;
		6'b111001: lut_value = 32'b10001010000101001101010101110101;
		6'b111010: lut_value = 32'b10001000100110000000111010000000;
		6'b111011: lut_value = 32'b10000111000111110110000110010110;
		6'b111100: lut_value = 32'b10000101101010101100001101100111;
		6'b111101: lut_value = 32'b10000100001110100010100011000011;
		6'b111110: lut_value = 32'b10000010110011011000011010011000;
		6'b111111: lut_value = 32'b10000001011001001101000111110011;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut2_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111101001110100100011011;
		6'b000010: lut_value = 32'b11111111111010011101001010110010;
		6'b000011: lut_value = 32'b11111111110111101011110011000100;
		6'b000100: lut_value = 32'b11111111110100111010011101010001;
		6'b000101: lut_value = 32'b11111111110010001001001001011001;
		6'b000110: lut_value = 32'b11111111101111010111110111011100;
		6'b000111: lut_value = 32'b11111111101100100110100111011001;
		6'b001000: lut_value = 32'b11111111101001110101011001010010;
		6'b001001: lut_value = 32'b11111111100111000100001101000101;
		6'b001010: lut_value = 32'b11111111100100010011000010110011;
		6'b001011: lut_value = 32'b11111111100001100001111010011100;
		6'b001100: lut_value = 32'b11111111011110110000110011111111;
		6'b001101: lut_value = 32'b11111111011011111111101111011110;
		6'b001110: lut_value = 32'b11111111011001001110101100110111;
		6'b001111: lut_value = 32'b11111111010110011101101100001010;
		6'b010000: lut_value = 32'b11111111010011101100101101011001;
		6'b010001: lut_value = 32'b11111111010000111011110000100010;
		6'b010010: lut_value = 32'b11111111001110001010110101100110;
		6'b010011: lut_value = 32'b11111111001011011001111100100100;
		6'b010100: lut_value = 32'b11111111001000101001000101011101;
		6'b010101: lut_value = 32'b11111111000101111000010000010001;
		6'b010110: lut_value = 32'b11111111000011000111011100111111;
		6'b010111: lut_value = 32'b11111111000000010110101011100111;
		6'b011000: lut_value = 32'b11111110111101100101111100001010;
		6'b011001: lut_value = 32'b11111110111010110101001110101000;
		6'b011010: lut_value = 32'b11111110111000000100100011000000;
		6'b011011: lut_value = 32'b11111110110101010011111001010011;
		6'b011100: lut_value = 32'b11111110110010100011010001100000;
		6'b011101: lut_value = 32'b11111110101111110010101011100111;
		6'b011110: lut_value = 32'b11111110101101000010000111101001;
		6'b011111: lut_value = 32'b11111110101010010001100101100101;
		6'b100000: lut_value = 32'b11111110100111100001000101011100;
		6'b100001: lut_value = 32'b11111110100100110000100111001101;
		6'b100010: lut_value = 32'b11111110100010000000001010111000;
		6'b100011: lut_value = 32'b11111110011111001111110000011110;
		6'b100100: lut_value = 32'b11111110011100011111010111111101;
		6'b100101: lut_value = 32'b11111110011001101111000001010111;
		6'b100110: lut_value = 32'b11111110010110111110101100101100;
		6'b100111: lut_value = 32'b11111110010100001110011001111010;
		6'b101000: lut_value = 32'b11111110010001011110001001000011;
		6'b101001: lut_value = 32'b11111110001110101101111010000110;
		6'b101010: lut_value = 32'b11111110001011111101101101000010;
		6'b101011: lut_value = 32'b11111110001001001101100001111010;
		6'b101100: lut_value = 32'b11111110000110011101011000101011;
		6'b101101: lut_value = 32'b11111110000011101101010001010110;
		6'b101110: lut_value = 32'b11111110000000111101001011111011;
		6'b101111: lut_value = 32'b11111101111110001101001000011011;
		6'b110000: lut_value = 32'b11111101111011011101000110110100;
		6'b110001: lut_value = 32'b11111101111000101101000111000111;
		6'b110010: lut_value = 32'b11111101110101111101001001010101;
		6'b110011: lut_value = 32'b11111101110011001101001101011100;
		6'b110100: lut_value = 32'b11111101110000011101010011011101;
		6'b110101: lut_value = 32'b11111101101101101101011011011001;
		6'b110110: lut_value = 32'b11111101101010111101100101001110;
		6'b110111: lut_value = 32'b11111101101000001101110000111101;
		6'b111000: lut_value = 32'b11111101100101011101111110100110;
		6'b111001: lut_value = 32'b11111101100010101110001110001000;
		6'b111010: lut_value = 32'b11111101011111111110011111100101;
		6'b111011: lut_value = 32'b11111101011101001110110010111011;
		6'b111100: lut_value = 32'b11111101011010011111001000001011;
		6'b111101: lut_value = 32'b11111101010111101111011111010101;
		6'b111110: lut_value = 32'b11111101010100111111111000011000;
		6'b111111: lut_value = 32'b11111101010010010000010011010110;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut3_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111101001110100011;
		6'b000010: lut_value = 32'b11111111111111111010011101000111;
		6'b000011: lut_value = 32'b11111111111111110111101011101010;
		6'b000100: lut_value = 32'b11111111111111110100111010001110;
		6'b000101: lut_value = 32'b11111111111111110010001000110001;
		6'b000110: lut_value = 32'b11111111111111101111010111010101;
		6'b000111: lut_value = 32'b11111111111111101100100101111001;
		6'b001000: lut_value = 32'b11111111111111101001110100011100;
		6'b001001: lut_value = 32'b11111111111111100111000011000000;
		6'b001010: lut_value = 32'b11111111111111100100010001100100;
		6'b001011: lut_value = 32'b11111111111111100001100000001000;
		6'b001100: lut_value = 32'b11111111111111011110101110101011;
		6'b001101: lut_value = 32'b11111111111111011011111101001111;
		6'b001110: lut_value = 32'b11111111111111011001001011110011;
		6'b001111: lut_value = 32'b11111111111111010110011010010111;
		6'b010000: lut_value = 32'b11111111111111010011101000111011;
		6'b010001: lut_value = 32'b11111111111111010000110111011111;
		6'b010010: lut_value = 32'b11111111111111001110000110000011;
		6'b010011: lut_value = 32'b11111111111111001011010100100111;
		6'b010100: lut_value = 32'b11111111111111001000100011001011;
		6'b010101: lut_value = 32'b11111111111111000101110001101111;
		6'b010110: lut_value = 32'b11111111111111000011000000010011;
		6'b010111: lut_value = 32'b11111111111111000000001110110111;
		6'b011000: lut_value = 32'b11111111111110111101011101011100;
		6'b011001: lut_value = 32'b11111111111110111010101100000000;
		6'b011010: lut_value = 32'b11111111111110110111111010100100;
		6'b011011: lut_value = 32'b11111111111110110101001001001000;
		6'b011100: lut_value = 32'b11111111111110110010010111101101;
		6'b011101: lut_value = 32'b11111111111110101111100110010001;
		6'b011110: lut_value = 32'b11111111111110101100110100110101;
		6'b011111: lut_value = 32'b11111111111110101010000011011010;
		6'b100000: lut_value = 32'b11111111111110100111010001111110;
		6'b100001: lut_value = 32'b11111111111110100100100000100011;
		6'b100010: lut_value = 32'b11111111111110100001101111000111;
		6'b100011: lut_value = 32'b11111111111110011110111101101100;
		6'b100100: lut_value = 32'b11111111111110011100001100010000;
		6'b100101: lut_value = 32'b11111111111110011001011010110101;
		6'b100110: lut_value = 32'b11111111111110010110101001011001;
		6'b100111: lut_value = 32'b11111111111110010011110111111110;
		6'b101000: lut_value = 32'b11111111111110010001000110100011;
		6'b101001: lut_value = 32'b11111111111110001110010101000111;
		6'b101010: lut_value = 32'b11111111111110001011100011101100;
		6'b101011: lut_value = 32'b11111111111110001000110010010001;
		6'b101100: lut_value = 32'b11111111111110000110000000110110;
		6'b101101: lut_value = 32'b11111111111110000011001111011010;
		6'b101110: lut_value = 32'b11111111111110000000011101111111;
		6'b101111: lut_value = 32'b11111111111101111101101100100100;
		6'b110000: lut_value = 32'b11111111111101111010111011001001;
		6'b110001: lut_value = 32'b11111111111101111000001001101110;
		6'b110010: lut_value = 32'b11111111111101110101011000010011;
		6'b110011: lut_value = 32'b11111111111101110010100110111000;
		6'b110100: lut_value = 32'b11111111111101101111110101011101;
		6'b110101: lut_value = 32'b11111111111101101101000100000010;
		6'b110110: lut_value = 32'b11111111111101101010010010100111;
		6'b110111: lut_value = 32'b11111111111101100111100001001100;
		6'b111000: lut_value = 32'b11111111111101100100101111110001;
		6'b111001: lut_value = 32'b11111111111101100001111110010110;
		6'b111010: lut_value = 32'b11111111111101011111001100111100;
		6'b111011: lut_value = 32'b11111111111101011100011011100001;
		6'b111100: lut_value = 32'b11111111111101011001101010000110;
		6'b111101: lut_value = 32'b11111111111101010110111000101011;
		6'b111110: lut_value = 32'b11111111111101010100000111010001;
		6'b111111: lut_value = 32'b11111111111101010001010101110110;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut4_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111111111101001110;
		6'b000010: lut_value = 32'b11111111111111111111111010011101;
		6'b000011: lut_value = 32'b11111111111111111111110111101011;
		6'b000100: lut_value = 32'b11111111111111111111110100111010;
		6'b000101: lut_value = 32'b11111111111111111111110010001000;
		6'b000110: lut_value = 32'b11111111111111111111101111010111;
		6'b000111: lut_value = 32'b11111111111111111111101100100101;
		6'b001000: lut_value = 32'b11111111111111111111101001110100;
		6'b001001: lut_value = 32'b11111111111111111111100111000010;
		6'b001010: lut_value = 32'b11111111111111111111100100010001;
		6'b001011: lut_value = 32'b11111111111111111111100001100000;
		6'b001100: lut_value = 32'b11111111111111111111011110101110;
		6'b001101: lut_value = 32'b11111111111111111111011011111101;
		6'b001110: lut_value = 32'b11111111111111111111011001001011;
		6'b001111: lut_value = 32'b11111111111111111111010110011010;
		6'b010000: lut_value = 32'b11111111111111111111010011101000;
		6'b010001: lut_value = 32'b11111111111111111111010000110111;
		6'b010010: lut_value = 32'b11111111111111111111001110000101;
		6'b010011: lut_value = 32'b11111111111111111111001011010100;
		6'b010100: lut_value = 32'b11111111111111111111001000100011;
		6'b010101: lut_value = 32'b11111111111111111111000101110001;
		6'b010110: lut_value = 32'b11111111111111111111000011000000;
		6'b010111: lut_value = 32'b11111111111111111111000000001110;
		6'b011000: lut_value = 32'b11111111111111111110111101011101;
		6'b011001: lut_value = 32'b11111111111111111110111010101011;
		6'b011010: lut_value = 32'b11111111111111111110110111111010;
		6'b011011: lut_value = 32'b11111111111111111110110101001000;
		6'b011100: lut_value = 32'b11111111111111111110110010010111;
		6'b011101: lut_value = 32'b11111111111111111110101111100110;
		6'b011110: lut_value = 32'b11111111111111111110101100110100;
		6'b011111: lut_value = 32'b11111111111111111110101010000011;
		6'b100000: lut_value = 32'b11111111111111111110100111010001;
		6'b100001: lut_value = 32'b11111111111111111110100100100000;
		6'b100010: lut_value = 32'b11111111111111111110100001101110;
		6'b100011: lut_value = 32'b11111111111111111110011110111101;
		6'b100100: lut_value = 32'b11111111111111111110011100001011;
		6'b100101: lut_value = 32'b11111111111111111110011001011010;
		6'b100110: lut_value = 32'b11111111111111111110010110101001;
		6'b100111: lut_value = 32'b11111111111111111110010011110111;
		6'b101000: lut_value = 32'b11111111111111111110010001000110;
		6'b101001: lut_value = 32'b11111111111111111110001110010100;
		6'b101010: lut_value = 32'b11111111111111111110001011100011;
		6'b101011: lut_value = 32'b11111111111111111110001000110001;
		6'b101100: lut_value = 32'b11111111111111111110000110000000;
		6'b101101: lut_value = 32'b11111111111111111110000011001110;
		6'b101110: lut_value = 32'b11111111111111111110000000011101;
		6'b101111: lut_value = 32'b11111111111111111101111101101100;
		6'b110000: lut_value = 32'b11111111111111111101111010111010;
		6'b110001: lut_value = 32'b11111111111111111101111000001001;
		6'b110010: lut_value = 32'b11111111111111111101110101010111;
		6'b110011: lut_value = 32'b11111111111111111101110010100110;
		6'b110100: lut_value = 32'b11111111111111111101101111110100;
		6'b110101: lut_value = 32'b11111111111111111101101101000011;
		6'b110110: lut_value = 32'b11111111111111111101101010010001;
		6'b110111: lut_value = 32'b11111111111111111101100111100000;
		6'b111000: lut_value = 32'b11111111111111111101100100101111;
		6'b111001: lut_value = 32'b11111111111111111101100001111101;
		6'b111010: lut_value = 32'b11111111111111111101011111001100;
		6'b111011: lut_value = 32'b11111111111111111101011100011010;
		6'b111100: lut_value = 32'b11111111111111111101011001101001;
		6'b111101: lut_value = 32'b11111111111111111101010110110111;
		6'b111110: lut_value = 32'b11111111111111111101010100000110;
		6'b111111: lut_value = 32'b11111111111111111101010001010100;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut5_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111111111111111101;
		6'b000010: lut_value = 32'b11111111111111111111111111111010;
		6'b000011: lut_value = 32'b11111111111111111111111111110111;
		6'b000100: lut_value = 32'b11111111111111111111111111110100;
		6'b000101: lut_value = 32'b11111111111111111111111111110010;
		6'b000110: lut_value = 32'b11111111111111111111111111101111;
		6'b000111: lut_value = 32'b11111111111111111111111111101100;
		6'b001000: lut_value = 32'b11111111111111111111111111101001;
		6'b001001: lut_value = 32'b11111111111111111111111111100111;
		6'b001010: lut_value = 32'b11111111111111111111111111100100;
		6'b001011: lut_value = 32'b11111111111111111111111111100001;
		6'b001100: lut_value = 32'b11111111111111111111111111011110;
		6'b001101: lut_value = 32'b11111111111111111111111111011011;
		6'b001110: lut_value = 32'b11111111111111111111111111011001;
		6'b001111: lut_value = 32'b11111111111111111111111111010110;
		6'b010000: lut_value = 32'b11111111111111111111111111010011;
		6'b010001: lut_value = 32'b11111111111111111111111111010000;
		6'b010010: lut_value = 32'b11111111111111111111111111001110;
		6'b010011: lut_value = 32'b11111111111111111111111111001011;
		6'b010100: lut_value = 32'b11111111111111111111111111001000;
		6'b010101: lut_value = 32'b11111111111111111111111111000101;
		6'b010110: lut_value = 32'b11111111111111111111111111000011;
		6'b010111: lut_value = 32'b11111111111111111111111111000000;
		6'b011000: lut_value = 32'b11111111111111111111111110111101;
		6'b011001: lut_value = 32'b11111111111111111111111110111010;
		6'b011010: lut_value = 32'b11111111111111111111111110110111;
		6'b011011: lut_value = 32'b11111111111111111111111110110101;
		6'b011100: lut_value = 32'b11111111111111111111111110110010;
		6'b011101: lut_value = 32'b11111111111111111111111110101111;
		6'b011110: lut_value = 32'b11111111111111111111111110101100;
		6'b011111: lut_value = 32'b11111111111111111111111110101010;
		6'b100000: lut_value = 32'b11111111111111111111111110100111;
		6'b100001: lut_value = 32'b11111111111111111111111110100100;
		6'b100010: lut_value = 32'b11111111111111111111111110100001;
		6'b100011: lut_value = 32'b11111111111111111111111110011110;
		6'b100100: lut_value = 32'b11111111111111111111111110011100;
		6'b100101: lut_value = 32'b11111111111111111111111110011001;
		6'b100110: lut_value = 32'b11111111111111111111111110010110;
		6'b100111: lut_value = 32'b11111111111111111111111110010011;
		6'b101000: lut_value = 32'b11111111111111111111111110010001;
		6'b101001: lut_value = 32'b11111111111111111111111110001110;
		6'b101010: lut_value = 32'b11111111111111111111111110001011;
		6'b101011: lut_value = 32'b11111111111111111111111110001000;
		6'b101100: lut_value = 32'b11111111111111111111111110000110;
		6'b101101: lut_value = 32'b11111111111111111111111110000011;
		6'b101110: lut_value = 32'b11111111111111111111111110000000;
		6'b101111: lut_value = 32'b11111111111111111111111101111101;
		6'b110000: lut_value = 32'b11111111111111111111111101111010;
		6'b110001: lut_value = 32'b11111111111111111111111101111000;
		6'b110010: lut_value = 32'b11111111111111111111111101110101;
		6'b110011: lut_value = 32'b11111111111111111111111101110010;
		6'b110100: lut_value = 32'b11111111111111111111111101101111;
		6'b110101: lut_value = 32'b11111111111111111111111101101101;
		6'b110110: lut_value = 32'b11111111111111111111111101101010;
		6'b110111: lut_value = 32'b11111111111111111111111101100111;
		6'b111000: lut_value = 32'b11111111111111111111111101100100;
		6'b111001: lut_value = 32'b11111111111111111111111101100001;
		6'b111010: lut_value = 32'b11111111111111111111111101011111;
		6'b111011: lut_value = 32'b11111111111111111111111101011100;
		6'b111100: lut_value = 32'b11111111111111111111111101011001;
		6'b111101: lut_value = 32'b11111111111111111111111101010110;
		6'b111110: lut_value = 32'b11111111111111111111111101010100;
		6'b111111: lut_value = 32'b11111111111111111111111101010001;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut6_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111111111111111111;
		6'b000010: lut_value = 32'b11111111111111111111111111111111;
		6'b000011: lut_value = 32'b11111111111111111111111111111111;
		6'b000100: lut_value = 32'b11111111111111111111111111111111;
		6'b000101: lut_value = 32'b11111111111111111111111111111111;
		6'b000110: lut_value = 32'b11111111111111111111111111111111;
		6'b000111: lut_value = 32'b11111111111111111111111111111111;
		6'b001000: lut_value = 32'b11111111111111111111111111111111;
		6'b001001: lut_value = 32'b11111111111111111111111111111111;
		6'b001010: lut_value = 32'b11111111111111111111111111111111;
		6'b001011: lut_value = 32'b11111111111111111111111111111111;
		6'b001100: lut_value = 32'b11111111111111111111111111111111;
		6'b001101: lut_value = 32'b11111111111111111111111111111111;
		6'b001110: lut_value = 32'b11111111111111111111111111111111;
		6'b001111: lut_value = 32'b11111111111111111111111111111111;
		6'b010000: lut_value = 32'b11111111111111111111111111111111;
		6'b010001: lut_value = 32'b11111111111111111111111111111111;
		6'b010010: lut_value = 32'b11111111111111111111111111111111;
		6'b010011: lut_value = 32'b11111111111111111111111111111111;
		6'b010100: lut_value = 32'b11111111111111111111111111111111;
		6'b010101: lut_value = 32'b11111111111111111111111111111111;
		6'b010110: lut_value = 32'b11111111111111111111111111111111;
		6'b010111: lut_value = 32'b11111111111111111111111111111111;
		6'b011000: lut_value = 32'b11111111111111111111111111111110;
		6'b011001: lut_value = 32'b11111111111111111111111111111110;
		6'b011010: lut_value = 32'b11111111111111111111111111111110;
		6'b011011: lut_value = 32'b11111111111111111111111111111110;
		6'b011100: lut_value = 32'b11111111111111111111111111111110;
		6'b011101: lut_value = 32'b11111111111111111111111111111110;
		6'b011110: lut_value = 32'b11111111111111111111111111111110;
		6'b011111: lut_value = 32'b11111111111111111111111111111110;
		6'b100000: lut_value = 32'b11111111111111111111111111111110;
		6'b100001: lut_value = 32'b11111111111111111111111111111110;
		6'b100010: lut_value = 32'b11111111111111111111111111111110;
		6'b100011: lut_value = 32'b11111111111111111111111111111110;
		6'b100100: lut_value = 32'b11111111111111111111111111111110;
		6'b100101: lut_value = 32'b11111111111111111111111111111110;
		6'b100110: lut_value = 32'b11111111111111111111111111111110;
		6'b100111: lut_value = 32'b11111111111111111111111111111110;
		6'b101000: lut_value = 32'b11111111111111111111111111111110;
		6'b101001: lut_value = 32'b11111111111111111111111111111110;
		6'b101010: lut_value = 32'b11111111111111111111111111111110;
		6'b101011: lut_value = 32'b11111111111111111111111111111110;
		6'b101100: lut_value = 32'b11111111111111111111111111111110;
		6'b101101: lut_value = 32'b11111111111111111111111111111110;
		6'b101110: lut_value = 32'b11111111111111111111111111111110;
		6'b101111: lut_value = 32'b11111111111111111111111111111101;
		6'b110000: lut_value = 32'b11111111111111111111111111111101;
		6'b110001: lut_value = 32'b11111111111111111111111111111101;
		6'b110010: lut_value = 32'b11111111111111111111111111111101;
		6'b110011: lut_value = 32'b11111111111111111111111111111101;
		6'b110100: lut_value = 32'b11111111111111111111111111111101;
		6'b110101: lut_value = 32'b11111111111111111111111111111101;
		6'b110110: lut_value = 32'b11111111111111111111111111111101;
		6'b110111: lut_value = 32'b11111111111111111111111111111101;
		6'b111000: lut_value = 32'b11111111111111111111111111111101;
		6'b111001: lut_value = 32'b11111111111111111111111111111101;
		6'b111010: lut_value = 32'b11111111111111111111111111111101;
		6'b111011: lut_value = 32'b11111111111111111111111111111101;
		6'b111100: lut_value = 32'b11111111111111111111111111111101;
		6'b111101: lut_value = 32'b11111111111111111111111111111101;
		6'b111110: lut_value = 32'b11111111111111111111111111111101;
		6'b111111: lut_value = 32'b11111111111111111111111111111101;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut7_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111111111111111111;
		6'b000010: lut_value = 32'b11111111111111111111111111111111;
		6'b000011: lut_value = 32'b11111111111111111111111111111111;
		6'b000100: lut_value = 32'b11111111111111111111111111111111;
		6'b000101: lut_value = 32'b11111111111111111111111111111111;
		6'b000110: lut_value = 32'b11111111111111111111111111111111;
		6'b000111: lut_value = 32'b11111111111111111111111111111111;
		6'b001000: lut_value = 32'b11111111111111111111111111111111;
		6'b001001: lut_value = 32'b11111111111111111111111111111111;
		6'b001010: lut_value = 32'b11111111111111111111111111111111;
		6'b001011: lut_value = 32'b11111111111111111111111111111111;
		6'b001100: lut_value = 32'b11111111111111111111111111111111;
		6'b001101: lut_value = 32'b11111111111111111111111111111111;
		6'b001110: lut_value = 32'b11111111111111111111111111111111;
		6'b001111: lut_value = 32'b11111111111111111111111111111111;
		6'b010000: lut_value = 32'b11111111111111111111111111111111;
		6'b010001: lut_value = 32'b11111111111111111111111111111111;
		6'b010010: lut_value = 32'b11111111111111111111111111111111;
		6'b010011: lut_value = 32'b11111111111111111111111111111111;
		6'b010100: lut_value = 32'b11111111111111111111111111111111;
		6'b010101: lut_value = 32'b11111111111111111111111111111111;
		6'b010110: lut_value = 32'b11111111111111111111111111111111;
		6'b010111: lut_value = 32'b11111111111111111111111111111111;
		6'b011000: lut_value = 32'b11111111111111111111111111111111;
		6'b011001: lut_value = 32'b11111111111111111111111111111111;
		6'b011010: lut_value = 32'b11111111111111111111111111111111;
		6'b011011: lut_value = 32'b11111111111111111111111111111111;
		6'b011100: lut_value = 32'b11111111111111111111111111111111;
		6'b011101: lut_value = 32'b11111111111111111111111111111111;
		6'b011110: lut_value = 32'b11111111111111111111111111111111;
		6'b011111: lut_value = 32'b11111111111111111111111111111111;
		6'b100000: lut_value = 32'b11111111111111111111111111111111;
		6'b100001: lut_value = 32'b11111111111111111111111111111111;
		6'b100010: lut_value = 32'b11111111111111111111111111111111;
		6'b100011: lut_value = 32'b11111111111111111111111111111111;
		6'b100100: lut_value = 32'b11111111111111111111111111111111;
		6'b100101: lut_value = 32'b11111111111111111111111111111111;
		6'b100110: lut_value = 32'b11111111111111111111111111111111;
		6'b100111: lut_value = 32'b11111111111111111111111111111111;
		6'b101000: lut_value = 32'b11111111111111111111111111111111;
		6'b101001: lut_value = 32'b11111111111111111111111111111111;
		6'b101010: lut_value = 32'b11111111111111111111111111111111;
		6'b101011: lut_value = 32'b11111111111111111111111111111111;
		6'b101100: lut_value = 32'b11111111111111111111111111111111;
		6'b101101: lut_value = 32'b11111111111111111111111111111111;
		6'b101110: lut_value = 32'b11111111111111111111111111111111;
		6'b101111: lut_value = 32'b11111111111111111111111111111111;
		6'b110000: lut_value = 32'b11111111111111111111111111111111;
		6'b110001: lut_value = 32'b11111111111111111111111111111111;
		6'b110010: lut_value = 32'b11111111111111111111111111111111;
		6'b110011: lut_value = 32'b11111111111111111111111111111111;
		6'b110100: lut_value = 32'b11111111111111111111111111111111;
		6'b110101: lut_value = 32'b11111111111111111111111111111111;
		6'b110110: lut_value = 32'b11111111111111111111111111111111;
		6'b110111: lut_value = 32'b11111111111111111111111111111111;
		6'b111000: lut_value = 32'b11111111111111111111111111111111;
		6'b111001: lut_value = 32'b11111111111111111111111111111111;
		6'b111010: lut_value = 32'b11111111111111111111111111111111;
		6'b111011: lut_value = 32'b11111111111111111111111111111111;
		6'b111100: lut_value = 32'b11111111111111111111111111111111;
		6'b111101: lut_value = 32'b11111111111111111111111111111111;
		6'b111110: lut_value = 32'b11111111111111111111111111111111;
		6'b111111: lut_value = 32'b11111111111111111111111111111111;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module Lut8_EXP
(
	input  wire [5:0]  index,
	output reg [31:0] lut_value
);

always @(*) begin
    case (index)
		6'b000000: lut_value = 32'b10000000000000000000000000000000;
		6'b000001: lut_value = 32'b11111111111111111111111111111111;
		6'b000010: lut_value = 32'b11111111111111111111111111111111;
		6'b000011: lut_value = 32'b11111111111111111111111111111111;
		6'b000100: lut_value = 32'b11111111111111111111111111111111;
		6'b000101: lut_value = 32'b11111111111111111111111111111111;
		6'b000110: lut_value = 32'b11111111111111111111111111111111;
		6'b000111: lut_value = 32'b11111111111111111111111111111111;
		6'b001000: lut_value = 32'b11111111111111111111111111111111;
		6'b001001: lut_value = 32'b11111111111111111111111111111111;
		6'b001010: lut_value = 32'b11111111111111111111111111111111;
		6'b001011: lut_value = 32'b11111111111111111111111111111111;
		6'b001100: lut_value = 32'b11111111111111111111111111111111;
		6'b001101: lut_value = 32'b11111111111111111111111111111111;
		6'b001110: lut_value = 32'b11111111111111111111111111111111;
		6'b001111: lut_value = 32'b11111111111111111111111111111111;
		6'b010000: lut_value = 32'b11111111111111111111111111111111;
		6'b010001: lut_value = 32'b11111111111111111111111111111111;
		6'b010010: lut_value = 32'b11111111111111111111111111111111;
		6'b010011: lut_value = 32'b11111111111111111111111111111111;
		6'b010100: lut_value = 32'b11111111111111111111111111111111;
		6'b010101: lut_value = 32'b11111111111111111111111111111111;
		6'b010110: lut_value = 32'b11111111111111111111111111111111;
		6'b010111: lut_value = 32'b11111111111111111111111111111111;
		6'b011000: lut_value = 32'b11111111111111111111111111111111;
		6'b011001: lut_value = 32'b11111111111111111111111111111111;
		6'b011010: lut_value = 32'b11111111111111111111111111111111;
		6'b011011: lut_value = 32'b11111111111111111111111111111111;
		6'b011100: lut_value = 32'b11111111111111111111111111111111;
		6'b011101: lut_value = 32'b11111111111111111111111111111111;
		6'b011110: lut_value = 32'b11111111111111111111111111111111;
		6'b011111: lut_value = 32'b11111111111111111111111111111111;
		6'b100000: lut_value = 32'b11111111111111111111111111111111;
		6'b100001: lut_value = 32'b11111111111111111111111111111111;
		6'b100010: lut_value = 32'b11111111111111111111111111111111;
		6'b100011: lut_value = 32'b11111111111111111111111111111111;
		6'b100100: lut_value = 32'b11111111111111111111111111111111;
		6'b100101: lut_value = 32'b11111111111111111111111111111111;
		6'b100110: lut_value = 32'b11111111111111111111111111111111;
		6'b100111: lut_value = 32'b11111111111111111111111111111111;
		6'b101000: lut_value = 32'b11111111111111111111111111111111;
		6'b101001: lut_value = 32'b11111111111111111111111111111111;
		6'b101010: lut_value = 32'b11111111111111111111111111111111;
		6'b101011: lut_value = 32'b11111111111111111111111111111111;
		6'b101100: lut_value = 32'b11111111111111111111111111111111;
		6'b101101: lut_value = 32'b11111111111111111111111111111111;
		6'b101110: lut_value = 32'b11111111111111111111111111111111;
		6'b101111: lut_value = 32'b11111111111111111111111111111111;
		6'b110000: lut_value = 32'b11111111111111111111111111111111;
		6'b110001: lut_value = 32'b11111111111111111111111111111111;
		6'b110010: lut_value = 32'b11111111111111111111111111111111;
		6'b110011: lut_value = 32'b11111111111111111111111111111111;
		6'b110100: lut_value = 32'b11111111111111111111111111111111;
		6'b110101: lut_value = 32'b11111111111111111111111111111111;
		6'b110110: lut_value = 32'b11111111111111111111111111111111;
		6'b110111: lut_value = 32'b11111111111111111111111111111111;
		6'b111000: lut_value = 32'b11111111111111111111111111111111;
		6'b111001: lut_value = 32'b11111111111111111111111111111111;
		6'b111010: lut_value = 32'b11111111111111111111111111111111;
		6'b111011: lut_value = 32'b11111111111111111111111111111111;
		6'b111100: lut_value = 32'b11111111111111111111111111111111;
		6'b111101: lut_value = 32'b11111111111111111111111111111111;
		6'b111110: lut_value = 32'b11111111111111111111111111111111;
		6'b111111: lut_value = 32'b11111111111111111111111111111111;
		default: lut_value = 32'd0;
    endcase
end
endmodule

module math_expf32(
	input wire clk,
	input wire rst_n,
	input wire iexp2_op_en,
	input wire [31:0] iexp2_rb,
	output wire iexp2_ra_en,
	output wire [31:0] iexp2_ra,
	output wire iexp2_luf_flag
);

reg exp_flag1, exp_flag2, exp_flag3, exp_flag4;
always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		exp_flag1 <= 1'b0;
		exp_flag2 <= 1'b0;
		exp_flag3 <= 1'b0;
		exp_flag4 <= 1'b0;
	end
	else begin
		exp_flag1 <= iexp2_op_en;
		exp_flag2 <= exp_flag1;
		exp_flag3 <= exp_flag2;
		exp_flag4 <= exp_flag3;
	end 
end 
    
wire [4:0] n;
wire [55:0] data_in;
wire [55:0] index;

assign data_in = {7'd0,1'b1,iexp2_rb[22:0],25'd0};
assign n = iexp2_rb[30]? (iexp2_rb[27:23]+1'b1) : (~iexp2_rb[27:23]);
assign index = iexp2_rb[30]? (data_in << n) : (data_in >> n);


reg over_flag, under_flag;
reg over_flag1  ;
reg under_flag1;
reg [31:0] reg_iexp2_rb;


reg [55:0] index_temp1, index_temp2;
always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		index_temp1 <= 56'd0;
	end 
	else if(iexp2_op_en)begin
		index_temp1 <= index;
	end
end 


always @(posedge clk or negedge rst_n) begin
  if(!rst_n) begin
    index_temp2 <= 1'd0;
  end
  else if(exp_flag1) begin
    index_temp2 <= index_temp1;
  end 
end

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		reg_iexp2_rb <= 32'd0;
	end
	else if(iexp2_op_en)begin
		reg_iexp2_rb <= iexp2_rb;
	end
end 

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		under_flag <= 1'b0;
	end
	else if(exp_flag1 && reg_iexp2_rb[30:23] > 8'd133 ) begin
		under_flag <= 1'b1;
	end
	else if(exp_flag1 && index_temp1[55:48] == 8'd127) begin
		under_flag <= 1'b1;
	end
	else if(exp_flag1 && index_temp1[55:48] == 8'd126 && index_temp1[47:0] != 48'd0) begin
		under_flag <= 1'b1;
	end 
	else begin
		under_flag <= 1'b0;
	end
end

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		over_flag <= 1'b0;
	end
	else if(exp_flag1 && reg_iexp2_rb[30:23] < 8'd102) begin
		over_flag <= 1'b1;
	end
	else begin
		over_flag <= 1'b0;
	end
end 

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		under_flag1 <= 1'b0;
	end
	else if(exp_flag2) begin
		under_flag1 <= under_flag;
	end
	else begin
		under_flag1 <= 1'd0;
	end 
end 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
  
always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		over_flag1 <= 1'b0;
	end
	else if(exp_flag2) begin
		over_flag1 <= over_flag;
	end
	else begin
		over_flag1 <= 1'b0;
	end 
end 

//cycle four
reg [7:0] reg_exp;
always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		reg_exp <= 8'd0;
	end 
	else if(exp_flag2 && index_temp2[55:48] < 8'd127 && index_temp2[47:0] == 48'd0) begin
		reg_exp <= 8'd127 - index_temp2[55:48];
	end 
	else if(exp_flag2 &&  index_temp2[55:48] < 8'd126) begin
		reg_exp <= 8'd126 - index_temp2[55:48];
	end 
	else begin
		reg_exp <= 8'd0;
	end 
end


wire [31:0] lut_A, lut_B, lut_C, lut_D, lut_E, lut_F, lut_G, lut_H;

Lut1_EXP Lut1_EXP
(
	.index		(index[47:42]),
	.lut_value	(lut_A)
);

Lut2_EXP Lut2_EXP
(
	.index		(index[41:36]),
	.lut_value 	(lut_B)
);

Lut3_EXP Lut3_EXP
(
	.index		(index[35:30]),
	.lut_value	(lut_C)
);

Lut4_EXP Lut4_EXP
(
	.index		(index[29:24]),
	.lut_value	(lut_D)
);

Lut5_EXP Lut5_EXP
(
	.index		(index[23:18]),
	.lut_value	(lut_E)
);

Lut6_EXP Lut6_EXP
(
	.index		(index[17:12]),
	.lut_value	(lut_F)
);

Lut7_EXP Lut7_EXP
(
	.index		(index[11:6]),
	.lut_value	(lut_G)
);

Lut8_EXP Lut8_EXP
(
	.index		(index[5:0]),
	.lut_value	(lut_H)
);

reg [31:0] A_tail, B_tail, C_tail, D_tail, E_tail, F_tail, G_tail, H_tail;

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		A_tail <= 32'd0;
		B_tail <= 32'd0;
		C_tail <= 32'd0;
		D_tail <= 32'd0;
		E_tail <= 32'd0;
		F_tail <= 32'd0;
		G_tail <= 32'd0;
		H_tail <= 32'd0;
	end
	else begin
		A_tail <= lut_A;
		B_tail <= lut_B;
		C_tail <= lut_C;
		D_tail <= lut_D;
		E_tail <= lut_E;
		F_tail <= lut_F;
		G_tail <= lut_G;
		H_tail <= lut_H;
	end 
end
 

wire [31:0] T1_tail, T2_tail, T3_tail, T4_tail;
reg [31:0] Rtail_T1, Rtail_T2, Rtail_T3, Rtail_T4;


mult_exp mult_one(
	.mult_a			(	A_tail		),
	.mult_b			(	B_tail		),
	.mult_c			(	T1_tail		)
);

mult_exp mult_two(
	.mult_a			(	C_tail		),
	.mult_b			(	D_tail		),
	.mult_c			(	T2_tail		)
);

mult_exp mult_three(
	.mult_a			(	E_tail		),
	.mult_b			(	F_tail		),
	.mult_c			(	T3_tail		)
);

mult_exp mult_four(
	.mult_a			(	G_tail		),
	.mult_b			(	H_tail		),
	.mult_c			(	T4_tail		)
);


always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		Rtail_T1 <= 32'd0;
		Rtail_T2 <= 32'd0;
		Rtail_T3 <= 32'd0;
		Rtail_T4 <= 32'd0;
	end 
	else begin
		Rtail_T1 <= T1_tail;
		Rtail_T2 <= T2_tail;
		Rtail_T3 <= T3_tail;
		Rtail_T4 <= T4_tail;
	end 
end 


wire [31:0] S1_tail, S2_tail;
reg [31:0] Rtail_S1, Rtail_S2;


mult_exp mult_five(
	.mult_a			(	Rtail_T1	),
	.mult_b			(	Rtail_T2	),
	.mult_c			(	S1_tail		)
);

mult_exp mult_six(
	.mult_a			(	Rtail_T3	),
	.mult_b			(	Rtail_T4	),
	.mult_c			(	S2_tail		)
);

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		Rtail_S1 <= 32'd0;
		Rtail_S2 <= 32'd0;
	end 
	else begin
		Rtail_S1 <= S1_tail;
		Rtail_S2 <= S2_tail;
	end 
end 

wire [31:0] Y_tail;

mult_exp mult_seven(
	.mult_a			(	Rtail_S1	),
	.mult_b			(	Rtail_S2	),
	.mult_c			(	Y_tail		)
);



reg [31:0] Result_exp;
always @(posedge clk or negedge rst_n) begin 
	if(!rst_n) begin
		Result_exp <= 32'd0;
	end 
	else if(under_flag1) begin
		Result_exp <= 32'd0;
	end
	else if(over_flag1) begin
		Result_exp <= 32'h3f800000;
	end
	else if(exp_flag3) begin
		Result_exp <= {1'd0, reg_exp, Y_tail[30:8]};
	end
	else begin
		Result_exp <= Result_exp;
	end 
end

assign iexp2_ra = Result_exp;
assign iexp2_ra_en = exp_flag4 ? 1'b1 : 1'b0;
assign iexp2_luf_flag = under_flag1? 1'b1 : 1'b0;
endmodule 